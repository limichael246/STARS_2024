`timescale 1ms/1ps

typedef enum logic [1:0] {
    INACTIVE = 2'b00,
    READY = 2'b01,
    ACTIVE = 2'b10
} VGA_state_t;

module tb;

    //Testbench parameters
    integer tb_test_num;
    string tb_test_case;

    

    // DUT Ports
    logic clk;
    logic nRst;

    //signals for controlling inputs/outputs
    logic mem_busy;
    VGA_state_t VGA_state;
    logic CPU_enable;

    //signals to/from VGA
    logic VGA_read;
    logic [31:0] VGA_adr;
    logic [31:0] data_to_VGA;

    //signals to/from UART
    logic UART_write;
    logic [31:0] UART_adr;
    logic [31:0] data_from_UART;

    //signals to/from CPU
    logic [31:0] CPU_instr_adr;
    logic [31:0] CPU_data_adr;
    logic CPU_read;
    logic CPU_write;
    logic [31:0] data_from_CPU;
    logic [3:0] CPU_sel;
    logic [31:0] instr_data_to_CPU;
    logic [31:0] data_to_CPU;

    //signals to/from memory/Wishbone
    logic [31:0] data_from_mem;
    logic mem_read;
    logic mem_write;
    logic [31:0] adr_to_mem;
    logic [31:0] data_to_mem;
    logic [3:0] sel_to_me;



    //Clock generation block
    localparam CLK_PERIOD = 10; // 100 Hz clk
    always begin
        clk = 1'b0;
        #(CLK_PERIOD / 2.0);
        clk = 1'b1;
        #(CLK_PERIOD / 2.0);
    end



    // DUT Instance
    request_handler2 reqhand (
        .clk(clk),
        .nRst(nRst),

        //signals for controlling inputs/outputs
        .mem_busy(mem_busy),
        .VGA_state(VGA_state),
        .CPU_enable(CPU_enable),

        //signals to/from VGA
        .VGA_read(VGA_read),
        .VGA_adr(VGA_adr),
        .data_to_VGA(data_to_VGA),

        //signals to/from UART
        .UART_write(UART_write),
        .UART_adr(UART_adr),
        .data_from_UART(data_to_UART),

        //signals to/from CPU
        .CPU_instr_adr(CPU_instr_adr),
        .CPU_data_adr(CPU_data_adr),
        .CPU_read(CPU_read),
        .CPU_write(CPU_write),
        .data_from_CPU(data_from_CPU),
        .CPU_sel(CPU_sel),
        .instr_data_to_CPU(instr_data_to_CPU),
        .data_to_CPU(data_to_CPU),

        //signals to/from memory/Wishbone
        .data_from_mem(data_from_mem),
        .mem_read(mem_read),
        .mem_write(mem_write),
        .adr_to_mem(adr_to_mem),
        .data_to_mem(data_to_mem),
        .sel_to_mem(sel_to_mem)
    );

    // Task to Check CPU_enable
    task check_;
        input logic expected_;
    begin
        if ( != ) begin
            $display("Error at test %d: %s", tb_test_num, tb_test_case);
            $display("Incorrect . Expected: %b, Actual: %b", , );
        end
    end
    endtask


    // Task to reset parameters
    task reset_parameters;
    begin
        nRst = 0;
        #10;
        nRst = 1;
        
    end
    endtask



    // Main test bench process
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, tb);

        


        $finish;
    end

endmodule
